module shape_rom(input  logic [4:0]  address,
					  output logic [15:0] shape
);

	parameter ADDR_WIDTH = 5;
	parameter DATA_WIDTH = 16;
	logic [ADDR_WIDTH-1:0] addr_reg;
	
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		//I
		16'b0100010001000100, 
		16'b0000000011110000, 
		16'b0010001000100010,
		16'b0000000011110000,
		//O
		16'b0000011001100000,
		16'b0000011001100000,
		16'b0000011001100000,
		16'b0000011001100000,
		//T
		16'b0000010011100000,
		16'b0000010001100100,
		16'b0000011100100000,
		16'b0000001001100010,
		//J
		16'b0000001000100110,
		16'b0000000001000111,
		16'b0000011001000100,
		16'b0000011100010000,
		//L
		16'b0000010001000110,
		16'b0000000001110100,
		16'b0000011000100010,
		16'b0000000001000111,
		//S
		16'b0000001101100000,
		16'b0100011000100000,
		16'b0000001101100000,
		16'b0100011000100000,
		//Z
		16'b0000110001100000,
		16'b0010011001000000,
		16'b0000110001100000,
		16'b0010011001000000
		};
		
	assign shape = ROM[address];
	
endmodule
